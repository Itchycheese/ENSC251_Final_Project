lib;
            Fand : out std_logic_vector(2 downto 0));
		Aand: in std_Logic;
Band: std_logic;

   F <= A ;
F;
Aand;
Fand;
Band;B;

